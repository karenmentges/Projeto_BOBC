module operativo (
    
);

endmodule